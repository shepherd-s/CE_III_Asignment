--Ejercicio 1.a (entity)
----------------------------

library ieee;
use ieee.std_logic_1164.all;

entity entity1 is
	port (f, g    : out std_logic;
	      x, y, z : in std_logic);
end entity entity1;
